/*
	Authored 2018-2019, Ryan Voo.

	All rights reserved.
	Redistribution and use in source and binary forms, with or without
	modification, are permitted provided that the following conditions
	are met:

	*	Redistributions of source code must retain the above
		copyright notice, this list of conditions and the following
		disclaimer.

	*	Redistributions in binary form must reproduce the above
		copyright notice, this list of conditions and the following
		disclaimer in the documentation and/or other materials
		provided with the distribution.

	*	Neither the name of the author nor the names of its
		contributors may be used to endorse or promote products
		derived from this software without specific prior written
		permission.

	THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
	"AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
	LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS
	FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
	COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,
	INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING,
	BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
	LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
	CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
	LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN
	ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
	POSSIBILITY OF SUCH DAMAGE.
*/

module data_mem(
	input			clk,
	input [31:0]		addr,
	input [31:0]		write_data,
	input			memwrite,
	input			memread,
	input [3:0]		sign_mask,
	output [31:0]		read_data,
	output reg [7:0]	led,
	output reg		clk_stall	/* Sets the clock high. */
);
	/*
	 *	Current state
	 */
	reg			state = 0;
	reg			operation_buf;

	/*
	 *	Possible states
	 */
	parameter		IDLE	= 0;
	parameter		OPERATE	= 1;

	parameter		READ	= 0;
	parameter		WRITE	= 1;


	/*
	 *	Line buffer
	 */
	reg [31:0]		word_buf;

	/*
	 *	Read buffer
	 */
	wire [31:0]		read_buf;

	/*
	 *	Buffers to store write data
	 */
	reg [31:0]		write_data_buffer;

	/*
	 *	Buffer to store address
	 */
	reg [31:0]		addr_buf;

	/*
	 *	Sign_mask buffer
	 */
	reg [3:0]		sign_mask_buf;

	/*
	 *	Block memory registers
	 *
	 *	(Bad practice: The constant for the size should be a `define).
	 */
	reg [31:0]		data_block[0:1023];

	/*
	 *	Wire assignments
	 */
	wire [9:0]		addr_block_addr;
	wire [9:0]		addr_buf_block_addr;
	wire [1:0]		addr_buf_byte_offset;

	wire [31:0]		replacement_word;

	/*
	 * Split the address into word index and byte index (within the selected
	 * word).
	 *
	 * BUG: The instruction memory supposedly occupies the first 0x1000
	 * addresses (hence the data memory starts at 0x1000), but we mask off
	 * the MSBs, so reads and writes to 0x100, 0x1100, and 0x2100 all end up
	 * at the same memory cell. This also implies that it's impossible to
	 * read/write to/from the instruction memory.
	 */
	assign			addr_block_addr		= addr[11:2];
	assign			addr_buf_block_addr	= addr_buf[11:2];
	assign			addr_buf_byte_offset	= addr_buf[1:0];

	/* Multiplexers. */
	reg			whole_word_read;

	mux2to1 read_mux(
		.input0(read_buf), /* Use combinatorial network output. */
		.input1(word_buf), /* Use memory output directly. */
		.select(whole_word_read),
		.out(read_data)
	);

	memory_multiplexer mem_mux(
		.addr_lsb(addr_buf_byte_offset),
		.word_buf(word_buf),
		.write_data_buffer(write_data_buffer),
		.sign_mask_buf(sign_mask_buf),
		.read_buf(read_buf),
		.replacement_word(replacement_word)
	);

	/*
	 *	This uses Yosys's support for nonzero initial values:
	 *
	 *		https://github.com/YosysHQ/yosys/commit/0793f1b196df536975a044a4ce53025c81d00c7f
	 *
	 *	Rather than using this simulation construct (`initial`),
	 *	the design should instead use a reset signal going to
	 *	modules in the design.
	 */
	initial begin
		$readmemh("verilog/data.hex", data_block);
		clk_stall = 0;
	end

	/*
	 *	LED register interfacing with I/O
	 */
	always @(posedge clk) begin
		if (memwrite == 1'b1 && addr == 32'h2000) begin
			led <= write_data[7:0];

			`ifdef SIMULATION_MODE
				/* Clock period is #2. */
				$display("@%0t cycles Writing to LED",
					$realtime / 2);
				if (write_data == 0) begin
					$writememh("memory_dump.hex", data_block);
					$finish;
				end
			`endif
		end
	end

	/*
	 *	State machine
	 */
	always @(posedge clk) begin
		case (state)
			IDLE: begin
				clk_stall <= 0;
				write_data_buffer <= write_data;
				addr_buf <= addr;
				sign_mask_buf <= sign_mask;

				word_buf <= data_block[addr_block_addr];

				if (memread == 1'b1) begin
					if (sign_mask[2:0] == 3'b111) begin
						whole_word_read <= 1'b1;
					end
					else begin
						whole_word_read <= 1'b0;
						clk_stall <= 1'b1;
						state <= OPERATE;
						operation_buf <= READ;
					end
				end
				else if (memwrite == 1'b1) begin
					clk_stall <= 1'b1;
					state <= OPERATE;
					operation_buf <= WRITE;
				end
			end

			OPERATE: begin
				if (operation_buf == WRITE)
					data_block[addr_buf_block_addr] <= replacement_word;

				clk_stall <= 1'b0;
				state <= IDLE;
			end
		endcase
	end
endmodule
